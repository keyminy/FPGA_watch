module hex2bcd_top(

);
reg st0,st1;
reg [4:0] cnt;
reg convert;


endmodule