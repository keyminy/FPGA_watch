module hex2bcd();

endmodule